class my_seq_item extends uvm_sequence_item;
`uvm_object_utils( my_seq_item )


function new();
  super.new;
endfunction


endclass
