interface my_if( input clk_i );

bit [3:0] cnt;

endinterface
