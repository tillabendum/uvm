package my_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"



`include "registers.sv"
`include "my_reg_file.sv"
`include "my_reg_block.sv"



`include "my_env.sv"
`include "my_test.sv"

endpackage
