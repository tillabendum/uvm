package my_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "my_obj.sv"
  `include "comp_a.sv"
  `include "comp_b.sv"
  `include "comp_c.sv"
  `include "comp_d.sv"
  `include "my_env.sv"
  `include "test.sv"

endpackage
