package my_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"


`include "comp_a.sv"
`include "comp_b.sv"
`include "comp_c.sv"
`include "my_env.sv"
`include "my_test.sv"

endpackage
