package my_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"


`include "my_seq_item.sv"
`include "my_sequence.sv"
`include "my_drv.sv"
`include "my_env.sv"
`include "my_test.sv"

endpackage
