package my_params_pkg;

localparam DWIDTH = 16;
localparam AWIDTH = 8;


endpackage
